class Generator;
    string name;

endclass